module scheduler #(
        parameter DATA_WIDTH = 64,
        parameter ADR_WIDTH =40,
        parameter HDR_WIDTH = 2
    )
    (
        ports
    );

endmodule
