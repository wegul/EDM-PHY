module sched (
    input wire [63:0] encoded_tx_data,
    input wire [1:0] encoded_tx_hdr,

    

);





endmodule