module test_eth_phy_tx;
    reg clk;
    reg [1:0] encoded_tx_hdr;
    reg [63:0] encoded_tx_data;

    


endmodule
